/home/shadab/shadab/libs/lefs/all.lef