

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO counter 
  PIN reset 
    ANTENNAPARTIALMETALAREA 3.024 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.448 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6696 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 10.7322 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 41.1272 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.403823 LAYER Via34 ;
  END reset
  PIN clk 
    ANTENNAPARTIALMETALAREA 11.9564 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.1666 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4824 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 34.2522 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 135.999 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 1.50222 LAYER Via23 ;
  END clk
  PIN count[7] 
    ANTENNADIFFAREA 0.56 LAYER Metal2 ; 
    ANTENNAPARTIALMETALAREA 3.346 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.667 LAYER Metal2 ;
  END count[7]
  PIN count[6] 
    ANTENNAPARTIALMETALAREA 4.942 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.709 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via23 ;
    ANTENNADIFFAREA 0.72 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.4376 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.328 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3924 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 15.0626 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 57.4766 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.74677 LAYER Via34 ;
  END count[6]
  PIN count[5] 
    ANTENNAPARTIALMETALAREA 6.659 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.592 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3924 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 24.4111 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 96.4976 LAYER Metal2 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via23 ;
    ANTENNAMAXCUTCAR 1.21793 LAYER Via23 ;
    ANTENNADIFFAREA 0.72 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.8784 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1936 LAYER Metal3 ;
    ANTENNAGATEAREA 0.3924 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 31.7465 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 125.024 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.21793 LAYER Via34 ;
  END count[5]
  PIN count[4] 
    ANTENNADIFFAREA 0.72 LAYER Metal2 ; 
    ANTENNAPARTIALMETALAREA 6.9612 LAYER Metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.9594 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3924 LAYER Metal2 ; 
    ANTENNAMAXAREACAR 23.3686 LAYER Metal2 ;
    ANTENNAMAXSIDEAREACAR 91.6283 LAYER Metal2 ;
    ANTENNAMAXCUTCAR 0.873385 LAYER Via23 ;
  END count[4]
  PIN count[3] 
    ANTENNADIFFAREA 0.72 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 4.7544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2956 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3924 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 49.5253 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 189.297 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.70707 LAYER Via34 ;
  END count[3]
  PIN count[2] 
    ANTENNADIFFAREA 0.72 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3924 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 45.1987 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 175.504 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.90702 LAYER Via56 ;
  END count[2]
  PIN count[1] 
    ANTENNADIFFAREA 0.72 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 9.1896 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.086 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2376 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 55.2685 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 210.439 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.70707 LAYER Via34 ;
  END count[1]
  PIN count[0] 
    ANTENNADIFFAREA 0.72 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4968 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 43.3305 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 165.589 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.68233 LAYER Via56 ;
  END count[0]
END counter

END LIBRARY
