/home/shadab/shadab/AdvGenusCUI_labs/MMMC/LEF/gsclib045_v3.5/lef/gsclib045_macro.lef